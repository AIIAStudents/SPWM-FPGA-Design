library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SPWM_index is
    generic (
        SIN_WIDTH      : integer := 9;     
        SIN_TABLE_SIZE : integer := 333
    );
    port(
        i_clk         : in  std_logic;       
        i_rst         : in  std_logic; 
        o_sin_value_a : out std_logic_vector(SIN_WIDTH-1 downto 0);
        o_sin_value_b : out std_logic_vector(SIN_WIDTH-1 downto 0);
        o_sin_value_c : out std_logic_vector(SIN_WIDTH-1 downto 0)
       --        o_sin_led     : out std_logic
    );
end entity;

architecture rtl of SPWM_index is
    -- 相位偏移量 = 0, 1/3 週期, 2/3 週期
    constant PHASE_A : integer := 0;
    constant PHASE_B : integer := SIN_TABLE_SIZE/3;
    constant PHASE_C : integer := 2*SIN_TABLE_SIZE/3;


    signal idx_a, idx_b, idx_c : std_logic_vector(SIN_WIDTH-1 downto 0);
    signal sin_index : unsigned(SIN_WIDTH-1 downto 0) := (others => '0');
    constant MAX_INDEX : unsigned(SIN_WIDTH-1 downto 0) := to_unsigned(SIN_TABLE_SIZE-1, SIN_WIDTH);


    type sine_table_type is array(0 to 332) of std_logic_vector(8 downto 0);
        constant sine_lut : sine_table_type := (
         0 => "001111111", 1 => "010000001", 2 => "010000100", 3 => "010000110",
         4 => "010001001", 5 => "010001011", 6 => "010001101", 7 => "010010000",
         8 => "010010010", 9 => "010010100", 10 => "010010111", 11 => "010011001",
         12 => "010011100", 13 => "010011110", 14 => "010100000", 15 => "010100010",
         16 => "010100101", 17 => "010100111", 18 => "010101001", 19 => "010101100",
         20 => "010101110", 21 => "010110000", 22 => "010110010", 23 => "010110100",
         24 => "010110111", 25 => "010111001", 26 => "010111011", 27 => "010111101",
         28 => "010111111", 29 => "011000001", 30 => "011000011", 31 => "011000101",
         32 => "011000111", 33 => "011001001", 34 => "011001011", 35 => "011001101",
         36 => "011001111", 37 => "011010001", 38 => "011010010", 39 => "011010100",
         40 => "011010110", 41 => "011011000", 42 => "011011001", 43 => "011011011",
         44 => "011011101", 45 => "011011110", 46 => "011100000", 47 => "011100001",
         48 => "011100011", 49 => "011100100", 50 => "011100110", 51 => "011100111",
         52 => "011101001", 53 => "011101010", 54 => "011101011", 55 => "011101100",
         56 => "011101110", 57 => "011101111", 58 => "011110000", 59 => "011110001",
         60 => "011110010", 61 => "011110011", 62 => "011110100", 63 => "011110101",
         64 => "011110110", 65 => "011110111", 66 => "011110111", 67 => "011111000",
         68 => "011111001", 69 => "011111001", 70 => "011111010", 71 => "011111011",
         72 => "011111011", 73 => "011111100", 74 => "011111100", 75 => "011111100",
         76 => "011111101", 77 => "011111101", 78 => "011111101", 79 => "011111110",
         80 => "011111110", 81 => "011111110", 82 => "011111110", 83 => "011111110",
         84 => "011111110", 85 => "011111110", 86 => "011111110", 87 => "011111110",
         88 => "011111101", 89 => "011111101", 90 => "011111101", 91 => "011111101",
         92 => "011111100", 93 => "011111100", 94 => "011111011", 95 => "011111011",
         96 => "011111010", 97 => "011111010", 98 => "011111001", 99 => "011111000",
         100 => "011111000", 101 => "011110111", 102 => "011110110", 103 => "011110101",
         104 => "011110100", 105 => "011110011", 106 => "011110010", 107 => "011110001",
         108 => "011110000", 109 => "011101111", 110 => "011101110", 111 => "011101101",
         112 => "011101100", 113 => "011101011", 114 => "011101001", 115 => "011101000",
         116 => "011100111", 117 => "011100101", 118 => "011100100", 119 => "011100010",
         120 => "011100001", 121 => "011011111", 122 => "011011110", 123 => "011011100",
         124 => "011011010", 125 => "011011001", 126 => "011010111", 127 => "011010101",
         128 => "011010011", 129 => "011010010", 130 => "011010000", 131 => "011001110",
         132 => "011001100", 133 => "011001010", 134 => "011001000", 135 => "011000110",
         136 => "011000100", 137 => "011000010", 138 => "011000000", 139 => "010111110",
         140 => "010111100", 141 => "010111010", 142 => "010111000", 143 => "010110101",
         144 => "010110011", 145 => "010110001", 146 => "010101111", 147 => "010101101",
         148 => "010101010", 149 => "010101000", 150 => "010100110", 151 => "010100100",
         152 => "010100001", 153 => "010011111", 154 => "010011101", 155 => "010011010",
         156 => "010011000", 157 => "010010110", 158 => "010010011", 159 => "010010001",
         160 => "010001111", 161 => "010001100", 162 => "010001010", 163 => "010000111",
         164 => "010000101", 165 => "010000011", 166 => "010000000", 167 => "001111110",
         168 => "001111011", 169 => "001111001", 170 => "001110111", 171 => "001110100",
         172 => "001110010", 173 => "001101111", 174 => "001101101", 175 => "001101011",
         176 => "001101000", 177 => "001100110", 178 => "001100100", 179 => "001100001",
         180 => "001011111", 181 => "001011101", 182 => "001011010", 183 => "001011000",
         184 => "001010110", 185 => "001010100", 186 => "001010001", 187 => "001001111",
         188 => "001001101", 189 => "001001011", 190 => "001001001", 191 => "001000110",
         192 => "001000100", 193 => "001000010", 194 => "001000000", 195 => "000111110",
         196 => "000111100", 197 => "000111010", 198 => "000111000", 199 => "000110110",
         200 => "000110100", 201 => "000110010", 202 => "000110000", 203 => "000101110",
         204 => "000101100", 205 => "000101011", 206 => "000101001", 207 => "000100111",
         208 => "000100101", 209 => "000100100", 210 => "000100010", 211 => "000100000",
         212 => "000011111", 213 => "000011101", 214 => "000011100", 215 => "000011010",
         216 => "000011001", 217 => "000010111", 218 => "000010110", 219 => "000010101",
         220 => "000010011", 221 => "000010010", 222 => "000010001", 223 => "000010000",
         224 => "000001111", 225 => "000001110", 226 => "000001101", 227 => "000001100",
         228 => "000001011", 229 => "000001010", 230 => "000001001", 231 => "000001000",
         232 => "000000111", 233 => "000000110", 234 => "000000110", 235 => "000000101",
         236 => "000000100", 237 => "000000100", 238 => "000000011", 239 => "000000011",
         240 => "000000010", 241 => "000000010", 242 => "000000001", 243 => "000000001",
         244 => "000000001", 245 => "000000001", 246 => "000000000", 247 => "000000000",
         248 => "000000000", 249 => "000000000", 250 => "000000000", 251 => "000000000",
         252 => "000000000", 253 => "000000000", 254 => "000000000", 255 => "000000001",
         256 => "000000001", 257 => "000000001", 258 => "000000010", 259 => "000000010",
         260 => "000000010", 261 => "000000011", 262 => "000000011", 263 => "000000100",
         264 => "000000101", 265 => "000000101", 266 => "000000110", 267 => "000000111",
         268 => "000000111", 269 => "000001000", 270 => "000001001", 271 => "000001010",
         272 => "000001011", 273 => "000001100", 274 => "000001101", 275 => "000001110",
         276 => "000001111", 277 => "000010000", 278 => "000010010", 279 => "000010011",
         280 => "000010100", 281 => "000010101", 282 => "000010111", 283 => "000011000",
         284 => "000011010", 285 => "000011011", 286 => "000011101", 287 => "000011110",
         288 => "000100000", 289 => "000100001", 290 => "000100011", 291 => "000100101",
         292 => "000100110", 293 => "000101000", 294 => "000101010", 295 => "000101100",
         296 => "000101101", 297 => "000101111", 298 => "000110001", 299 => "000110011",
         300 => "000110101", 301 => "000110111", 302 => "000111001", 303 => "000111011",
         304 => "000111101", 305 => "000111111", 306 => "001000001", 307 => "001000011",
         308 => "001000101", 309 => "001000111", 310 => "001001010", 311 => "001001100",
         312 => "001001110", 313 => "001010000", 314 => "001010010", 315 => "001010101",
         316 => "001010111", 317 => "001011001", 318 => "001011100", 319 => "001011110",
         320 => "001100000", 321 => "001100010", 322 => "001100101", 323 => "001100111",
         324 => "001101010", 325 => "001101100", 326 => "001101110", 327 => "001110001",
         328 => "001110011", 329 => "001110101", 330 => "001111000", 331 => "001111010",
         332 => "001111101"
);


begin

    phase_acc: process(i_clk, i_rst)
    begin
        if i_rst = '0' then
            sin_index <= (others => '0');
        elsif rising_edge(i_clk) then
            if sin_index = MAX_INDEX then
                sin_index <= (others => '0');
            else
                sin_index <= sin_index + 1;
            end if;
        end if;
    end process;

    idx_a <= std_logic_vector(to_unsigned( (to_integer(unsigned(sin_index)) + PHASE_A) mod SIN_TABLE_SIZE, SIN_WIDTH));
    idx_b <= std_logic_vector(to_unsigned( (to_integer(unsigned(sin_index)) + PHASE_B) mod SIN_TABLE_SIZE, SIN_WIDTH));
    idx_c <= std_logic_vector(to_unsigned( (to_integer(unsigned(sin_index)) + PHASE_C) mod SIN_TABLE_SIZE, SIN_WIDTH));



    o_sin_value_a <= sine_lut( to_integer(unsigned(idx_a)) );
    o_sin_value_b <= sine_lut( to_integer(unsigned(idx_b)) );
    o_sin_value_c <= sine_lut( to_integer(unsigned(idx_c)) );


--    sin_LED : process(sin_index)
--    begin
--        if sin_index < to_unsigned(SIN_TABLE_SIZE/2, SIN_WIDTH) then
--            o_sin_led <= '1';  
--        else
--            o_sin_led <= '0'; 
--        end if;
--    end process;';

end architecture;
