library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity SPWM_index is
    generic (
        SIN_WIDTH      : integer := 9;     
        SIN_TABLE_SIZE : integer := 333
    );
    port(
        i_clk         : in  std_logic;       
        i_rst         : in  std_logic; 
        o_sin_value_a : out std_logic_vector(7 downto 0);
        o_sin_value_b : out std_logic_vector(7 downto 0);
        o_sin_value_c : out std_logic_vector(7 downto 0)
       --        o_sin_led     : out std_logic
    );
end entity;

architecture rtl of SPWM_index is
    -- 相位偏移量 = 0, 1/3 週期, 2/3 週期
    constant PHASE_A : integer := 0;
    constant PHASE_B : integer := SIN_TABLE_SIZE/3;
    constant PHASE_C : integer := 2*SIN_TABLE_SIZE/3;

    signal idx_a, idx_b, idx_c : std_logic_vector(SIN_WIDTH-1 downto 0);
    signal sin_index           : std_logic_vector(SIN_WIDTH-1 downto 0) ;

    type sine_table_type is array(0 to 332) of std_logic_vector(7 downto 0);
    constant sine_lut : sine_table_type := (
        0 => "10000000", 1 => "10000010", 2 => "10000100", 3 => "10000111", 4 => "10001001",
        5 => "10001100", 6 => "10001110", 7 => "10010000", 8 => "10010011", 9 => "10010101",
        10 => "10010111", 11 => "10011010", 12 => "10011100", 13 => "10011110", 14 => "10100001",
        15 => "10100011", 16 => "10100101", 17 => "10101000", 18 => "10101010", 19 => "10101100",
        20 => "10101110", 21 => "10110001", 22 => "10110011", 23 => "10110101", 24 => "10110111",
        25 => "10111001", 26 => "10111100", 27 => "10111110", 28 => "11000000", 29 => "11000010",
        30 => "11000100", 31 => "11000110", 32 => "11001000", 33 => "11001010", 34 => "11001100",
        35 => "11001110", 36 => "11010000", 37 => "11010001", 38 => "11010011", 39 => "11010101",
        40 => "11010111", 41 => "11011001", 42 => "11011010", 43 => "11011100", 44 => "11011110",
        45 => "11011111", 46 => "11100001", 47 => "11100010", 48 => "11100100", 49 => "11100101",
        50 => "11100111", 51 => "11101000", 52 => "11101001", 53 => "11101011", 54 => "11101100",
        55 => "11101101", 56 => "11101111", 57 => "11110000", 58 => "11110001", 59 => "11110010",
        60 => "11110011", 61 => "11110100", 62 => "11110101", 63 => "11110110", 64 => "11110111",
        65 => "11111000", 66 => "11111000", 67 => "11111001", 68 => "11111010", 69 => "11111010",
        70 => "11111011", 71 => "11111100", 72 => "11111100", 73 => "11111101", 74 => "11111101",
        75 => "11111101", 76 => "11111110", 77 => "11111110", 78 => "11111110", 79 => "11111111",
        80 => "11111111", 81 => "11111111", 82 => "11111111", 83 => "11111111", 84 => "11111111",
        85 => "11111111", 86 => "11111111", 87 => "11111111", 88 => "11111110", 89 => "11111110",
        90 => "11111110", 91 => "11111110", 92 => "11111101", 93 => "11111101", 94 => "11111100",
        95 => "11111100", 96 => "11111011", 97 => "11111011", 98 => "11111010", 99 => "11111001",
        100 => "11111001", 101 => "11111000", 102 => "11110111", 103 => "11110110", 104 => "11110101",
        105 => "11110100", 106 => "11110011", 107 => "11110010", 108 => "11110001", 109 => "11110000",
        110 => "11101111", 111 => "11101110", 112 => "11101101", 113 => "11101011", 114 => "11101010",
        115 => "11101001", 116 => "11100111", 117 => "11100110", 118 => "11100101", 119 => "11100011",
        120 => "11100010", 121 => "11100000", 122 => "11011110", 123 => "11011101", 124 => "11011011",
        125 => "11011001", 126 => "11011000", 127 => "11010110", 128 => "11010100", 129 => "11010010",
        130 => "11010001", 131 => "11001111", 132 => "11001101", 133 => "11001011", 134 => "11001001",
        135 => "11000111", 136 => "11000101", 137 => "11000011", 138 => "11000001", 139 => "10111111",
        140 => "10111101", 141 => "10111011", 142 => "10111000", 143 => "10110110", 144 => "10110100",
        145 => "10110010", 146 => "10110000", 147 => "10101101", 148 => "10101011", 149 => "10101001",
        150 => "10100111", 151 => "10100100", 152 => "10100010", 153 => "10100000", 154 => "10011101",
        155 => "10011011", 156 => "10011001", 157 => "10010110", 158 => "10010100", 159 => "10010001",
        160 => "10001111", 161 => "10001101", 162 => "10001010", 163 => "10001000", 164 => "10000110",
        165 => "10000011", 166 => "10000001", 167 => "01111110", 168 => "01111100", 169 => "01111001",
        170 => "01110111", 171 => "01110101", 172 => "01110010", 173 => "01110000", 174 => "01101110",
        175 => "01101011", 176 => "01101001", 177 => "01100110", 178 => "01100100", 179 => "01100010",
        180 => "01011111", 181 => "01011101", 182 => "01011011", 183 => "01011000", 184 => "01010110",
        185 => "01010100", 186 => "01010010", 187 => "01001111", 188 => "01001101", 189 => "01001011",
        190 => "01001001", 191 => "01000111", 192 => "01000100", 193 => "01000010", 194 => "01000000",
        195 => "00111110", 196 => "00111100", 197 => "00111010", 198 => "00111000", 199 => "00110110",
        200 => "00110100", 201 => "00110010", 202 => "00110000", 203 => "00101110", 204 => "00101101",
        205 => "00101011", 206 => "00101001", 207 => "00100111", 208 => "00100110", 209 => "00100100",
        210 => "00100010", 211 => "00100001", 212 => "00011111", 213 => "00011101", 214 => "00011100",
        215 => "00011010", 216 => "00011001", 217 => "00011000", 218 => "00010110", 219 => "00010101",
        220 => "00010100", 221 => "00010010", 222 => "00010001", 223 => "00010000", 224 => "00001111",
        225 => "00001110", 226 => "00001101", 227 => "00001100", 228 => "00001011", 229 => "00001010",
        230 => "00001001", 231 => "00001000", 232 => "00000111", 233 => "00000110", 234 => "00000110",
        235 => "00000101", 236 => "00000100", 237 => "00000100", 238 => "00000011", 239 => "00000011",
        240 => "00000010", 241 => "00000010", 242 => "00000001", 243 => "00000001", 244 => "00000001",
        245 => "00000001", 246 => "00000000", 247 => "00000000", 248 => "00000000", 249 => "00000000",
        250 => "00000000", 251 => "00000000", 252 => "00000000", 253 => "00000000", 254 => "00000000",
        255 => "00000001", 256 => "00000001", 257 => "00000001", 258 => "00000010", 259 => "00000010",
        260 => "00000010", 261 => "00000011", 262 => "00000011", 263 => "00000100", 264 => "00000101",
        265 => "00000101", 266 => "00000110", 267 => "00000111", 268 => "00000111", 269 => "00001000",
        270 => "00001001", 271 => "00001010", 272 => "00001011", 273 => "00001100", 274 => "00001101",
        275 => "00001110", 276 => "00001111", 277 => "00010000", 278 => "00010010", 279 => "00010011",
        280 => "00010100", 281 => "00010110", 282 => "00010111", 283 => "00011000", 284 => "00011010",
        285 => "00011011", 286 => "00011101", 287 => "00011110", 288 => "00100000", 289 => "00100001",
        290 => "00100011", 291 => "00100101", 292 => "00100110", 293 => "00101000", 294 => "00101010",
        295 => "00101100", 296 => "00101110", 297 => "00101111", 298 => "00110001", 299 => "00110011",
        300 => "00110101", 301 => "00110111", 302 => "00111001", 303 => "00111011", 304 => "00111101",
        305 => "00111111", 306 => "01000001", 307 => "01000011", 308 => "01000110", 309 => "01001000",
        310 => "01001010", 311 => "01001100", 312 => "01001110", 313 => "01010001", 314 => "01010011",
        315 => "01010101", 316 => "01010111", 317 => "01011010", 318 => "01011100", 319 => "01011110",
        320 => "01100001", 321 => "01100011", 322 => "01100101", 323 => "01101000", 324 => "01101010",
        325 => "01101100", 326 => "01101111", 327 => "01110001", 328 => "01110011", 329 => "01110110",
        330 => "01111000", 331 => "01111011", 332 => "01111101"
    );


begin

    phase_acc: process(i_clk, i_rst)
    begin
        if i_rst = '0' then
            sin_index <= (others => '0');
        elsif rising_edge(i_clk) then
            if sin_index = std_logic_vector(to_unsigned(SIN_TABLE_SIZE - 1, sin_index'length)) then
                sin_index <= (others => '0');
            else
                sin_index <= sin_index + "1";
            end if;
        end if;
    end process;

    idx_a <= sin_index;
    idx_b <= std_logic_vector(to_unsigned( (to_integer(unsigned(sin_index)) + PHASE_B) mod SIN_TABLE_SIZE, SIN_WIDTH));
    idx_c <= std_logic_vector(to_unsigned( (to_integer(unsigned(sin_index)) + PHASE_C) mod SIN_TABLE_SIZE, SIN_WIDTH));



    o_sin_value_a <= sine_lut( to_integer(unsigned(idx_a)) );
    o_sin_value_b <= sine_lut( to_integer(unsigned(idx_b)) );
    o_sin_value_c <= sine_lut( to_integer(unsigned(idx_c)) );

--    sin_LED : process(sin_index)
--    begin
--        if sin_index < to_unsigned(SIN_TABLE_SIZE/2, SIN_WIDTH) then
--            o_sin_led <= '1';  
--        else
--            o_sin_led <= '0'; 
--        end if;
--    end process;';

end architecture;
