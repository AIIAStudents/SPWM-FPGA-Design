library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SPWM_main is
    generic (
        SIN_WIDTH         : integer := 8;
      	SIN_TABLE_SIZE     : integer := 256;
        SIN_UPDATE_PERIOD : integer := 1
    );
    port(
        i_clk        : in  std_logic;
        i_rst        : in  std_logic;
        i_sw_freq   : in  std_logic_vector(3 downto 0); 
        o_pwm_out    : out std_logic;
        o_sin_led    : out std_logic
    );
end entity;

architecture rtl of SPWM_main is

    type STATE_TYPE is (STATE_HIGH, STATE_LOW);
    signal STATE : STATE_TYPE := STATE_LOW;
    signal step_val : unsigned(SIN_WIDTH-1 downto 0) := (others=>'0');
    signal sin_index  : unsigned(SIN_WIDTH-1 downto 0) := (others => '0');
    signal sin_value  : unsigned(SIN_WIDTH-1 downto 0);
    signal cnt_high   : integer range 0 to 2**SIN_WIDTH-1 := 0;
    signal cnt_low    : integer range 0 to 2**SIN_WIDTH-1 := 0;
    signal cnt_sin    : integer := 0;

    type sine_table_type is array(0 to 255) of unsigned(7 downto 0);
        constant sine_lut : sine_table_type := (
        0 => "01111111", 1 => "10000010", 2 => "10000101", 3 => "10001000",
        4 => "10001011", 5 => "10001111", 6 => "10010010", 7 => "10010101",
        8 => "10011000", 9 => "10011011", 10 => "10011110", 11 => "10100001",
        12 => "10100100", 13 => "10100111", 14 => "10101010", 15 => "10101101",
        16 => "10110000", 17 => "10110011", 18 => "10110110", 19 => "10111000",
        20 => "10111011", 21 => "10111110", 22 => "11000001", 23 => "11000011",
        24 => "11000110", 25 => "11001000", 26 => "11001011", 27 => "11001101",
        28 => "11010000", 29 => "11010010", 30 => "11010101", 31 => "11010111",
        32 => "11011001", 33 => "11011011", 34 => "11011101", 35 => "11100000",
        36 => "11100010", 37 => "11100100", 38 => "11100101", 39 => "11100111",
        40 => "11101001", 41 => "11101011", 42 => "11101100", 43 => "11101110",
        44 => "11101111", 45 => "11110001", 46 => "11110010", 47 => "11110100",
        48 => "11110101", 49 => "11110110", 50 => "11110111", 51 => "11111000",
        52 => "11111001", 53 => "11111010", 54 => "11111011", 55 => "11111011",
        56 => "11111100", 57 => "11111101", 58 => "11111101", 59 => "11111110",
        60 => "11111110", 61 => "11111110", 62 => "11111110", 63 => "11111110",
        64 => "11111111", 65 => "11111110", 66 => "11111110", 67 => "11111110",
        68 => "11111110", 69 => "11111110", 70 => "11111101", 71 => "11111101",
        72 => "11111100", 73 => "11111011", 74 => "11111011", 75 => "11111010",
        76 => "11111001", 77 => "11111000", 78 => "11110111", 79 => "11110110",
        80 => "11110101", 81 => "11110100", 82 => "11110010", 83 => "11110001",
        84 => "11101111", 85 => "11101110", 86 => "11101100", 87 => "11101011",
        88 => "11101001", 89 => "11100111", 90 => "11100101", 91 => "11100100",
        92 => "11100010", 93 => "11100000", 94 => "11011101", 95 => "11011011",
        96 => "11011001", 97 => "11010111", 98 => "11010101", 99 => "11010010",
        100 => "11010000", 101 => "11001101", 102 => "11001011", 103 => "11001000",
        104 => "11000110", 105 => "11000011", 106 => "11000001", 107 => "10111110",
        108 => "10111011", 109 => "10111000", 110 => "10110110", 111 => "10110011",
        112 => "10110000", 113 => "10101101", 114 => "10101010", 115 => "10100111",
        116 => "10100100", 117 => "10100001", 118 => "10011110", 119 => "10011011",
        120 => "10011000", 121 => "10010101", 122 => "10010010", 123 => "10001111",
        124 => "10001011", 125 => "10001000", 126 => "10000101", 127 => "10000010",
        128 => "01111111", 129 => "01111100", 130 => "01111001", 131 => "01110110",
        132 => "01110011", 133 => "01101111", 134 => "01101100", 135 => "01101001",
        136 => "01100110", 137 => "01100011", 138 => "01100000", 139 => "01011101",
        140 => "01011010", 141 => "01010111", 142 => "01010100", 143 => "01010001",
        144 => "01001110", 145 => "01001011", 146 => "01001000", 147 => "01000110",
        148 => "01000011", 149 => "01000000", 150 => "00111101", 151 => "00111011",
        152 => "00111000", 153 => "00110110", 154 => "00110011", 155 => "00110001",
        156 => "00101110", 157 => "00101100", 158 => "00101001", 159 => "00100111",
        160 => "00100101", 161 => "00100011", 162 => "00100001", 163 => "00011110",
        164 => "00011100", 165 => "00011010", 166 => "00011001", 167 => "00010111",
        168 => "00010101", 169 => "00010011", 170 => "00010010", 171 => "00010000",
        172 => "00001111", 173 => "00001101", 174 => "00001100", 175 => "00001010",
        176 => "00001001", 177 => "00001000", 178 => "00000111", 179 => "00000110",
        180 => "00000101", 181 => "00000100", 182 => "00000011", 183 => "00000011",
        184 => "00000010", 185 => "00000001", 186 => "00000001", 187 => "00000000",
        188 => "00000000", 189 => "00000000", 190 => "00000000", 191 => "00000000",
        192 => "00000000", 193 => "00000000", 194 => "00000000", 195 => "00000000",
        196 => "00000000", 197 => "00000000", 198 => "00000001", 199 => "00000001",
        200 => "00000010", 201 => "00000011", 202 => "00000011", 203 => "00000100",
        204 => "00000101", 205 => "00000110", 206 => "00000111", 207 => "00001000",
        208 => "00001001", 209 => "00001010", 210 => "00001100", 211 => "00001101",
        212 => "00001111", 213 => "00010000", 214 => "00010010", 215 => "00010011",
        216 => "00010101", 217 => "00010111", 218 => "00011001", 219 => "00011010",
        220 => "00011100", 221 => "00011110", 222 => "00100001", 223 => "00100011",
        224 => "00100101", 225 => "00100111", 226 => "00101001", 227 => "00101100",
        228 => "00101110", 229 => "00110001", 230 => "00110011", 231 => "00110110",
        232 => "00111000", 233 => "00111011", 234 => "00111101", 235 => "01000000",
        236 => "01000011", 237 => "01000110", 238 => "01001000", 239 => "01001011",
        240 => "01001110", 241 => "01010001", 242 => "01010100", 243 => "01010111",
        244 => "01011010", 245 => "01011101", 246 => "01100000", 247 => "01100011",
        248 => "01100110", 249 => "01101001", 250 => "01101100", 251 => "01101111",
        252 => "01110011", 253 => "01110110", 254 => "01111001", 255 => "01111100"
    );


begin

    lut_proc : process(sin_index)
    begin
        sin_value <= sine_lut(to_integer(sin_index));
    end process;
    
    sin_LED : process(sin_index)
    begin
        if sin_index < to_unsigned(SIN_TABLE_SIZE/2, SIN_WIDTH) then
            o_sin_led <= '1';  
        else
            o_sin_led <= '0'; 
        end if;
    end process;
    
  process(i_sw_freq)
  begin
    step_val <= to_unsigned(2 ** to_integer(unsigned(i_sw_freq)), SIN_WIDTH);
  end process;

    counter_high : process(i_clk, i_rst)
    begin 
        if (i_rst = '0') then
            cnt_high <= 0;
        elsif rising_edge(i_clk) then
            if (STATE = STATE_HIGH) then
                if  (cnt_high < ((to_integer(sin_value)))) then
                    cnt_high <= cnt_high + 1;
                else
                    cnt_high <= 0;
                end if;
            else
                cnt_high <= 0;
            end if;
        end if;
    end process;

    counter_low : process(i_clk, i_rst)
    begin
        if (i_rst = '0') then
            cnt_low <= 0;
        elsif rising_edge(i_clk) then
            if (STATE = STATE_LOW) then
                if (cnt_low < (((2**SIN_WIDTH - 1 - to_integer(sin_value))))) then
                    cnt_low <= cnt_low + 1;
                else
                    cnt_low <= 0;
                end if;
            else
                cnt_low <= 0;
            end if;
        end if;
    end process;

    fsm_proc : process(i_clk, i_rst)
    begin
        if (i_rst = '0') then
            STATE     <= STATE_LOW;
            sin_index <= (others => '0');
            cnt_sin   <= 0;
        elsif rising_edge(i_clk) then
            case STATE is
                when STATE_HIGH =>
                    if (cnt_high = ((to_integer(sin_value) ))) then
                        STATE <= STATE_LOW;
                    end if;

                when STATE_LOW =>
                    if (cnt_low = ((2**SIN_WIDTH - 1 - to_integer(sin_value)))) then 
                        STATE <= STATE_HIGH;
                        if (cnt_sin = SIN_UPDATE_PERIOD - 1) then
                            cnt_sin <= 0;
                            if (sin_index = to_unsigned(SIN_TABLE_SIZE-1, SIN_WIDTH)) then
                                sin_index <= (others => '0');
                            else
                               sin_index <= sin_index  + step_val;
                            end if;
                        else
                            cnt_sin <= cnt_sin + 1;
                        end if;
                    end if;
            end case;
        end if;
    end process;


    outt : process(state)
    begin
        if (state = STATE_HIGH) then
            o_pwm_out <= '1';
        else
            o_pwm_out <= '0';
        end if;
    end process;

end architecture;
